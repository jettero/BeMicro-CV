// bemicro_cv.v

// Generated using ACDS version 14.0 200 at 2014.10.29.21:49:07

`timescale 1 ps / 1 ps
module bemicro_cv (
		output wire [7:0]  led_export,                    //         led.export
		input  wire [2:0]  sw_export,                     //          sw.export
		input  wire [1:0]  pb_export,                     //          pb.export
		output wire [12:0] ddr3_mem_a,                    //        ddr3.mem_a
		output wire [2:0]  ddr3_mem_ba,                   //            .mem_ba
		output wire [0:0]  ddr3_mem_ck,                   //            .mem_ck
		output wire [0:0]  ddr3_mem_ck_n,                 //            .mem_ck_n
		output wire [0:0]  ddr3_mem_cke,                  //            .mem_cke
		output wire [0:0]  ddr3_mem_cs_n,                 //            .mem_cs_n
		output wire [1:0]  ddr3_mem_dm,                   //            .mem_dm
		output wire [0:0]  ddr3_mem_ras_n,                //            .mem_ras_n
		output wire [0:0]  ddr3_mem_cas_n,                //            .mem_cas_n
		output wire [0:0]  ddr3_mem_we_n,                 //            .mem_we_n
		output wire        ddr3_mem_reset_n,              //            .mem_reset_n
		inout  wire [15:0] ddr3_mem_dq,                   //            .mem_dq
		inout  wire [1:0]  ddr3_mem_dqs,                  //            .mem_dqs
		inout  wire [1:0]  ddr3_mem_dqs_n,                //            .mem_dqs_n
		output wire [0:0]  ddr3_mem_odt,                  //            .mem_odt
		input  wire        reset_reset_n,                 //       reset.reset_n
		input  wire        ddr3_oct_rzqin,                //    ddr3_oct.rzqin
		output wire        ddr3_status_local_init_done,   // ddr3_status.local_init_done
		output wire        ddr3_status_local_cal_success, //            .local_cal_success
		output wire        ddr3_status_local_cal_fail,    //            .local_cal_fail
		input  wire        clk_clk                        //         clk.clk
	);

	wire         syspll_outclk0_clk;                                        // syspll:outclk_0 -> [LED:clk, ddr3_control:mp_cmd_clk_0_clk, ddr3_control:mp_rfifo_clk_0_clk, ddr3_control:mp_wfifo_clk_0_clk, dip_sw:clk, irq_mapper:clk, jtag_uart:clk, mm_bridge_0:clk, mm_interconnect_0:syspll_outclk0_clk, mm_interconnect_1:syspll_outclk0_clk, nios_cpu:clk, onchip_mem:clk, pb_sw:clk, rst_controller:clk, sys_clk_timer:clk, sysid:clock]
	wire   [3:0] nios_cpu_instruction_master_burstcount;                    // nios_cpu:i_burstcount -> mm_interconnect_0:nios_cpu_instruction_master_burstcount
	wire         nios_cpu_instruction_master_waitrequest;                   // mm_interconnect_0:nios_cpu_instruction_master_waitrequest -> nios_cpu:i_waitrequest
	wire  [27:0] nios_cpu_instruction_master_address;                       // nios_cpu:i_address -> mm_interconnect_0:nios_cpu_instruction_master_address
	wire         nios_cpu_instruction_master_read;                          // nios_cpu:i_read -> mm_interconnect_0:nios_cpu_instruction_master_read
	wire  [31:0] nios_cpu_instruction_master_readdata;                      // mm_interconnect_0:nios_cpu_instruction_master_readdata -> nios_cpu:i_readdata
	wire         nios_cpu_instruction_master_readdatavalid;                 // mm_interconnect_0:nios_cpu_instruction_master_readdatavalid -> nios_cpu:i_readdatavalid
	wire   [3:0] nios_cpu_data_master_burstcount;                           // nios_cpu:d_burstcount -> mm_interconnect_0:nios_cpu_data_master_burstcount
	wire         nios_cpu_data_master_waitrequest;                          // mm_interconnect_0:nios_cpu_data_master_waitrequest -> nios_cpu:d_waitrequest
	wire  [31:0] nios_cpu_data_master_writedata;                            // nios_cpu:d_writedata -> mm_interconnect_0:nios_cpu_data_master_writedata
	wire  [27:0] nios_cpu_data_master_address;                              // nios_cpu:d_address -> mm_interconnect_0:nios_cpu_data_master_address
	wire         nios_cpu_data_master_write;                                // nios_cpu:d_write -> mm_interconnect_0:nios_cpu_data_master_write
	wire         nios_cpu_data_master_read;                                 // nios_cpu:d_read -> mm_interconnect_0:nios_cpu_data_master_read
	wire  [31:0] nios_cpu_data_master_readdata;                             // mm_interconnect_0:nios_cpu_data_master_readdata -> nios_cpu:d_readdata
	wire         nios_cpu_data_master_debugaccess;                          // nios_cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios_cpu_data_master_debugaccess
	wire         nios_cpu_data_master_readdatavalid;                        // mm_interconnect_0:nios_cpu_data_master_readdatavalid -> nios_cpu:d_readdatavalid
	wire   [3:0] nios_cpu_data_master_byteenable;                           // nios_cpu:d_byteenable -> mm_interconnect_0:nios_cpu_data_master_byteenable
	wire         mm_interconnect_0_nios_cpu_jtag_debug_module_waitrequest;  // nios_cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:nios_cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios_cpu_jtag_debug_module_writedata;    // mm_interconnect_0:nios_cpu_jtag_debug_module_writedata -> nios_cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios_cpu_jtag_debug_module_address;      // mm_interconnect_0:nios_cpu_jtag_debug_module_address -> nios_cpu:jtag_debug_module_address
	wire         mm_interconnect_0_nios_cpu_jtag_debug_module_write;        // mm_interconnect_0:nios_cpu_jtag_debug_module_write -> nios_cpu:jtag_debug_module_write
	wire         mm_interconnect_0_nios_cpu_jtag_debug_module_read;         // mm_interconnect_0:nios_cpu_jtag_debug_module_read -> nios_cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios_cpu_jtag_debug_module_readdata;     // nios_cpu:jtag_debug_module_readdata -> mm_interconnect_0:nios_cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios_cpu_jtag_debug_module_debugaccess;  // mm_interconnect_0:nios_cpu_jtag_debug_module_debugaccess -> nios_cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios_cpu_jtag_debug_module_byteenable;   // mm_interconnect_0:nios_cpu_jtag_debug_module_byteenable -> nios_cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_writedata;                 // mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire  [13:0] mm_interconnect_0_onchip_mem_s1_address;                   // mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	wire         mm_interconnect_0_onchip_mem_s1_chipselect;                // mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire         mm_interconnect_0_onchip_mem_s1_clken;                     // mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	wire         mm_interconnect_0_onchip_mem_s1_write;                     // mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_readdata;                  // onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_mem_s1_byteenable;                // mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         mm_interconnect_0_ddr3_control_avl_0_waitrequest;          // ddr3_control:avl_ready_0 -> mm_interconnect_0:ddr3_control_avl_0_waitrequest
	wire   [2:0] mm_interconnect_0_ddr3_control_avl_0_burstcount;           // mm_interconnect_0:ddr3_control_avl_0_burstcount -> ddr3_control:avl_size_0
	wire  [31:0] mm_interconnect_0_ddr3_control_avl_0_writedata;            // mm_interconnect_0:ddr3_control_avl_0_writedata -> ddr3_control:avl_wdata_0
	wire  [24:0] mm_interconnect_0_ddr3_control_avl_0_address;              // mm_interconnect_0:ddr3_control_avl_0_address -> ddr3_control:avl_addr_0
	wire         mm_interconnect_0_ddr3_control_avl_0_write;                // mm_interconnect_0:ddr3_control_avl_0_write -> ddr3_control:avl_write_req_0
	wire         mm_interconnect_0_ddr3_control_avl_0_beginbursttransfer;   // mm_interconnect_0:ddr3_control_avl_0_beginbursttransfer -> ddr3_control:avl_burstbegin_0
	wire         mm_interconnect_0_ddr3_control_avl_0_read;                 // mm_interconnect_0:ddr3_control_avl_0_read -> ddr3_control:avl_read_req_0
	wire  [31:0] mm_interconnect_0_ddr3_control_avl_0_readdata;             // ddr3_control:avl_rdata_0 -> mm_interconnect_0:ddr3_control_avl_0_readdata
	wire         mm_interconnect_0_ddr3_control_avl_0_readdatavalid;        // ddr3_control:avl_rdata_valid_0 -> mm_interconnect_0:ddr3_control_avl_0_readdatavalid
	wire   [3:0] mm_interconnect_0_ddr3_control_avl_0_byteenable;           // mm_interconnect_0:ddr3_control_avl_0_byteenable -> ddr3_control:avl_be_0
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;              // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;               // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [9:0] mm_interconnect_0_mm_bridge_0_s0_address;                  // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                    // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                     // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                 // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;              // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;            // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;               // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire   [0:0] mm_bridge_0_m0_burstcount;                                 // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire         mm_bridge_0_m0_waitrequest;                                // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [9:0] mm_bridge_0_m0_address;                                    // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire  [31:0] mm_bridge_0_m0_writedata;                                  // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                      // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire         mm_bridge_0_m0_read;                                       // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire  [31:0] mm_bridge_0_m0_readdata;                                   // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire   [3:0] mm_bridge_0_m0_byteenable;                                 // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                              // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;             // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                        // mm_interconnect_1:LED_s1_writedata -> LED:writedata
	wire   [1:0] mm_interconnect_1_led_s1_address;                          // mm_interconnect_1:LED_s1_address -> LED:address
	wire         mm_interconnect_1_led_s1_chipselect;                       // mm_interconnect_1:LED_s1_chipselect -> LED:chipselect
	wire         mm_interconnect_1_led_s1_write;                            // mm_interconnect_1:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                         // LED:readdata -> mm_interconnect_1:LED_s1_readdata
	wire   [1:0] mm_interconnect_1_pb_sw_s1_address;                        // mm_interconnect_1:pb_sw_s1_address -> pb_sw:address
	wire  [31:0] mm_interconnect_1_pb_sw_s1_readdata;                       // pb_sw:readdata -> mm_interconnect_1:pb_sw_s1_readdata
	wire   [1:0] mm_interconnect_1_dip_sw_s1_address;                       // mm_interconnect_1:dip_sw_s1_address -> dip_sw:address
	wire  [31:0] mm_interconnect_1_dip_sw_s1_readdata;                      // dip_sw:readdata -> mm_interconnect_1:dip_sw_s1_readdata
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;              // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;             // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                  // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;               // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire         irq_mapper_receiver0_irq;                                  // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_cpu_d_irq_irq;                                        // irq_mapper:sender_irq -> nios_cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [LED:reset_n, ddr3_control:mp_cmd_reset_n_0_reset_n, dip_sw:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_bridge_0:reset, mm_interconnect_0:nios_cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, nios_cpu:reset_n, onchip_mem:reset, pb_sw:reset_n, rst_translator:in_reset, sys_clk_timer:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios_cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [ddr3_control:global_reset_n, syspll:rst]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [ddr3_control:mp_rfifo_reset_n_0_reset_n, ddr3_control:mp_wfifo_reset_n_0_reset_n, ddr3_control:soft_reset_n, rst_controller:reset_in0]
	wire         nios_cpu_jtag_debug_module_reset_reset;                    // nios_cpu:jtag_debug_module_resetrequest -> rst_controller_002:reset_in1

	bemicro_cv_nios_cpu nios_cpu (
		.clk                                   (syspll_outclk0_clk),                                       //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (nios_cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios_cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios_cpu_data_master_read),                                //                          .read
		.d_readdata                            (nios_cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios_cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios_cpu_data_master_write),                               //                          .write
		.d_writedata                           (nios_cpu_data_master_writedata),                           //                          .writedata
		.d_burstcount                          (nios_cpu_data_master_burstcount),                          //                          .burstcount
		.d_readdatavalid                       (nios_cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios_cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios_cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (nios_cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios_cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_burstcount                          (nios_cpu_instruction_master_burstcount),                   //                          .burstcount
		.i_readdatavalid                       (nios_cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios_cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                          // custom_instruction_master.readra
	);

	bemicro_cv_onchip_mem onchip_mem (
		.clk        (syspll_outclk0_clk),                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	bemicro_cv_sys_clk_timer sys_clk_timer (
		.clk        (syspll_outclk0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	bemicro_cv_jtag_uart jtag_uart (
		.clk            (syspll_outclk0_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	bemicro_cv_sysid sysid (
		.clock    (syspll_outclk0_clk),                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	bemicro_cv_dip_sw dip_sw (
		.clk      (syspll_outclk0_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_dip_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_dip_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                             // external_connection.export
	);

	bemicro_cv_LED led (
		.clk        (syspll_outclk0_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	bemicro_cv_pb_sw pb_sw (
		.clk      (syspll_outclk0_clk),                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_1_pb_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pb_sw_s1_readdata), //                    .readdata
		.in_port  (pb_export)                            // external_connection.export
	);

	bemicro_cv_ddr3_control ddr3_control (
		.pll_ref_clk                (clk_clk),                                                 //        pll_ref_clk.clk
		.global_reset_n             (~rst_controller_001_reset_out_reset),                     //       global_reset.reset_n
		.soft_reset_n               (~rst_controller_002_reset_out_reset),                     //         soft_reset.reset_n
		.afi_clk                    (),                                                        //            afi_clk.clk
		.afi_half_clk               (),                                                        //       afi_half_clk.clk
		.afi_reset_n                (),                                                        //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                        //   afi_reset_export.reset_n
		.mem_a                      (ddr3_mem_a),                                              //             memory.mem_a
		.mem_ba                     (ddr3_mem_ba),                                             //                   .mem_ba
		.mem_ck                     (ddr3_mem_ck),                                             //                   .mem_ck
		.mem_ck_n                   (ddr3_mem_ck_n),                                           //                   .mem_ck_n
		.mem_cke                    (ddr3_mem_cke),                                            //                   .mem_cke
		.mem_cs_n                   (ddr3_mem_cs_n),                                           //                   .mem_cs_n
		.mem_dm                     (ddr3_mem_dm),                                             //                   .mem_dm
		.mem_ras_n                  (ddr3_mem_ras_n),                                          //                   .mem_ras_n
		.mem_cas_n                  (ddr3_mem_cas_n),                                          //                   .mem_cas_n
		.mem_we_n                   (ddr3_mem_we_n),                                           //                   .mem_we_n
		.mem_reset_n                (ddr3_mem_reset_n),                                        //                   .mem_reset_n
		.mem_dq                     (ddr3_mem_dq),                                             //                   .mem_dq
		.mem_dqs                    (ddr3_mem_dqs),                                            //                   .mem_dqs
		.mem_dqs_n                  (ddr3_mem_dqs_n),                                          //                   .mem_dqs_n
		.mem_odt                    (ddr3_mem_odt),                                            //                   .mem_odt
		.avl_ready_0                (mm_interconnect_0_ddr3_control_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_0_ddr3_control_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_0_ddr3_control_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_0_ddr3_control_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_0_ddr3_control_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_0_ddr3_control_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_0_ddr3_control_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_0_ddr3_control_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_0_ddr3_control_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_0_ddr3_control_avl_0_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (syspll_outclk0_clk),                                      //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (~rst_controller_reset_out_reset),                         //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (syspll_outclk0_clk),                                      //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (~rst_controller_002_reset_out_reset),                     // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (syspll_outclk0_clk),                                      //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (~rst_controller_002_reset_out_reset),                     // mp_wfifo_reset_n_0.reset_n
		.local_init_done            (ddr3_status_local_init_done),                             //             status.local_init_done
		.local_cal_success          (ddr3_status_local_cal_success),                           //                   .local_cal_success
		.local_cal_fail             (ddr3_status_local_cal_fail),                              //                   .local_cal_fail
		.oct_rzqin                  (ddr3_oct_rzqin),                                          //                oct.rzqin
		.pll_mem_clk                (),                                                        //        pll_sharing.pll_mem_clk
		.pll_write_clk              (),                                                        //                   .pll_write_clk
		.pll_locked                 (),                                                        //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (),                                                        //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (),                                                        //                   .pll_addr_cmd_clk
		.pll_avl_clk                (),                                                        //                   .pll_avl_clk
		.pll_config_clk             (),                                                        //                   .pll_config_clk
		.pll_dr_clk                 (),                                                        //                   .pll_dr_clk
		.pll_dr_clk_pre_phy_clk     (),                                                        //                   .pll_dr_clk_pre_phy_clk
		.pll_mem_phy_clk            (),                                                        //                   .pll_mem_phy_clk
		.afi_phy_clk                (),                                                        //                   .afi_phy_clk
		.pll_avl_phy_clk            ()                                                         //                   .pll_avl_phy_clk
	);

	bemicro_cv_syspll syspll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (syspll_outclk0_clk),                 // outclk0.clk
		.outclk_1 (),                                   // outclk1.clk
		.locked   ()                                    //  locked.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (syspll_outclk0_clk),                             //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)                      //      .debugaccess
	);

	bemicro_cv_mm_interconnect_0 mm_interconnect_0 (
		.syspll_outclk0_clk                           (syspll_outclk0_clk),                                       //                         syspll_outclk0.clk
		.nios_cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // nios_cpu_reset_n_reset_bridge_in_reset.reset
		.nios_cpu_data_master_address                 (nios_cpu_data_master_address),                             //                   nios_cpu_data_master.address
		.nios_cpu_data_master_waitrequest             (nios_cpu_data_master_waitrequest),                         //                                       .waitrequest
		.nios_cpu_data_master_burstcount              (nios_cpu_data_master_burstcount),                          //                                       .burstcount
		.nios_cpu_data_master_byteenable              (nios_cpu_data_master_byteenable),                          //                                       .byteenable
		.nios_cpu_data_master_read                    (nios_cpu_data_master_read),                                //                                       .read
		.nios_cpu_data_master_readdata                (nios_cpu_data_master_readdata),                            //                                       .readdata
		.nios_cpu_data_master_readdatavalid           (nios_cpu_data_master_readdatavalid),                       //                                       .readdatavalid
		.nios_cpu_data_master_write                   (nios_cpu_data_master_write),                               //                                       .write
		.nios_cpu_data_master_writedata               (nios_cpu_data_master_writedata),                           //                                       .writedata
		.nios_cpu_data_master_debugaccess             (nios_cpu_data_master_debugaccess),                         //                                       .debugaccess
		.nios_cpu_instruction_master_address          (nios_cpu_instruction_master_address),                      //            nios_cpu_instruction_master.address
		.nios_cpu_instruction_master_waitrequest      (nios_cpu_instruction_master_waitrequest),                  //                                       .waitrequest
		.nios_cpu_instruction_master_burstcount       (nios_cpu_instruction_master_burstcount),                   //                                       .burstcount
		.nios_cpu_instruction_master_read             (nios_cpu_instruction_master_read),                         //                                       .read
		.nios_cpu_instruction_master_readdata         (nios_cpu_instruction_master_readdata),                     //                                       .readdata
		.nios_cpu_instruction_master_readdatavalid    (nios_cpu_instruction_master_readdatavalid),                //                                       .readdatavalid
		.ddr3_control_avl_0_address                   (mm_interconnect_0_ddr3_control_avl_0_address),             //                     ddr3_control_avl_0.address
		.ddr3_control_avl_0_write                     (mm_interconnect_0_ddr3_control_avl_0_write),               //                                       .write
		.ddr3_control_avl_0_read                      (mm_interconnect_0_ddr3_control_avl_0_read),                //                                       .read
		.ddr3_control_avl_0_readdata                  (mm_interconnect_0_ddr3_control_avl_0_readdata),            //                                       .readdata
		.ddr3_control_avl_0_writedata                 (mm_interconnect_0_ddr3_control_avl_0_writedata),           //                                       .writedata
		.ddr3_control_avl_0_beginbursttransfer        (mm_interconnect_0_ddr3_control_avl_0_beginbursttransfer),  //                                       .beginbursttransfer
		.ddr3_control_avl_0_burstcount                (mm_interconnect_0_ddr3_control_avl_0_burstcount),          //                                       .burstcount
		.ddr3_control_avl_0_byteenable                (mm_interconnect_0_ddr3_control_avl_0_byteenable),          //                                       .byteenable
		.ddr3_control_avl_0_readdatavalid             (mm_interconnect_0_ddr3_control_avl_0_readdatavalid),       //                                       .readdatavalid
		.ddr3_control_avl_0_waitrequest               (~mm_interconnect_0_ddr3_control_avl_0_waitrequest),        //                                       .waitrequest
		.mm_bridge_0_s0_address                       (mm_interconnect_0_mm_bridge_0_s0_address),                 //                         mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                         (mm_interconnect_0_mm_bridge_0_s0_write),                   //                                       .write
		.mm_bridge_0_s0_read                          (mm_interconnect_0_mm_bridge_0_s0_read),                    //                                       .read
		.mm_bridge_0_s0_readdata                      (mm_interconnect_0_mm_bridge_0_s0_readdata),                //                                       .readdata
		.mm_bridge_0_s0_writedata                     (mm_interconnect_0_mm_bridge_0_s0_writedata),               //                                       .writedata
		.mm_bridge_0_s0_burstcount                    (mm_interconnect_0_mm_bridge_0_s0_burstcount),              //                                       .burstcount
		.mm_bridge_0_s0_byteenable                    (mm_interconnect_0_mm_bridge_0_s0_byteenable),              //                                       .byteenable
		.mm_bridge_0_s0_readdatavalid                 (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),           //                                       .readdatavalid
		.mm_bridge_0_s0_waitrequest                   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),             //                                       .waitrequest
		.mm_bridge_0_s0_debugaccess                   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),             //                                       .debugaccess
		.nios_cpu_jtag_debug_module_address           (mm_interconnect_0_nios_cpu_jtag_debug_module_address),     //             nios_cpu_jtag_debug_module.address
		.nios_cpu_jtag_debug_module_write             (mm_interconnect_0_nios_cpu_jtag_debug_module_write),       //                                       .write
		.nios_cpu_jtag_debug_module_read              (mm_interconnect_0_nios_cpu_jtag_debug_module_read),        //                                       .read
		.nios_cpu_jtag_debug_module_readdata          (mm_interconnect_0_nios_cpu_jtag_debug_module_readdata),    //                                       .readdata
		.nios_cpu_jtag_debug_module_writedata         (mm_interconnect_0_nios_cpu_jtag_debug_module_writedata),   //                                       .writedata
		.nios_cpu_jtag_debug_module_byteenable        (mm_interconnect_0_nios_cpu_jtag_debug_module_byteenable),  //                                       .byteenable
		.nios_cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_nios_cpu_jtag_debug_module_waitrequest), //                                       .waitrequest
		.nios_cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_nios_cpu_jtag_debug_module_debugaccess), //                                       .debugaccess
		.onchip_mem_s1_address                        (mm_interconnect_0_onchip_mem_s1_address),                  //                          onchip_mem_s1.address
		.onchip_mem_s1_write                          (mm_interconnect_0_onchip_mem_s1_write),                    //                                       .write
		.onchip_mem_s1_readdata                       (mm_interconnect_0_onchip_mem_s1_readdata),                 //                                       .readdata
		.onchip_mem_s1_writedata                      (mm_interconnect_0_onchip_mem_s1_writedata),                //                                       .writedata
		.onchip_mem_s1_byteenable                     (mm_interconnect_0_onchip_mem_s1_byteenable),               //                                       .byteenable
		.onchip_mem_s1_chipselect                     (mm_interconnect_0_onchip_mem_s1_chipselect),               //                                       .chipselect
		.onchip_mem_s1_clken                          (mm_interconnect_0_onchip_mem_s1_clken)                     //                                       .clken
	);

	bemicro_cv_mm_interconnect_1 mm_interconnect_1 (
		.syspll_outclk0_clk                            (syspll_outclk0_clk),                                        //                          syspll_outclk0.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                    //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                 //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                 //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                       //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                   //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                              //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                      //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                  //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                //                                        .debugaccess
		.dip_sw_s1_address                             (mm_interconnect_1_dip_sw_s1_address),                       //                               dip_sw_s1.address
		.dip_sw_s1_readdata                            (mm_interconnect_1_dip_sw_s1_readdata),                      //                                        .readdata
		.jtag_uart_avalon_jtag_slave_address           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_avalon_jtag_slave_read              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.LED_s1_address                                (mm_interconnect_1_led_s1_address),                          //                                  LED_s1.address
		.LED_s1_write                                  (mm_interconnect_1_led_s1_write),                            //                                        .write
		.LED_s1_readdata                               (mm_interconnect_1_led_s1_readdata),                         //                                        .readdata
		.LED_s1_writedata                              (mm_interconnect_1_led_s1_writedata),                        //                                        .writedata
		.LED_s1_chipselect                             (mm_interconnect_1_led_s1_chipselect),                       //                                        .chipselect
		.pb_sw_s1_address                              (mm_interconnect_1_pb_sw_s1_address),                        //                                pb_sw_s1.address
		.pb_sw_s1_readdata                             (mm_interconnect_1_pb_sw_s1_readdata),                       //                                        .readdata
		.sys_clk_timer_s1_address                      (mm_interconnect_1_sys_clk_timer_s1_address),                //                        sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                        (mm_interconnect_1_sys_clk_timer_s1_write),                  //                                        .write
		.sys_clk_timer_s1_readdata                     (mm_interconnect_1_sys_clk_timer_s1_readdata),               //                                        .readdata
		.sys_clk_timer_s1_writedata                    (mm_interconnect_1_sys_clk_timer_s1_writedata),              //                                        .writedata
		.sys_clk_timer_s1_chipselect                   (mm_interconnect_1_sys_clk_timer_s1_chipselect),             //                                        .chipselect
		.sysid_control_slave_address                   (mm_interconnect_1_sysid_control_slave_address),             //                     sysid_control_slave.address
		.sysid_control_slave_readdata                  (mm_interconnect_1_sysid_control_slave_readdata)             //                                        .readdata
	);

	bemicro_cv_irq_mapper irq_mapper (
		.clk           (syspll_outclk0_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_cpu_d_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (rst_controller_002_reset_out_reset), // reset_in0.reset
		.clk            (syspll_outclk0_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios_cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
